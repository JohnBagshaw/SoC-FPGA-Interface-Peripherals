module SPI_interface (sclk, clk, din, dout, data_out, clock_out, chipsel);
